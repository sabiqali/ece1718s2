module mv_gen(input [7:0] c, input [7:0] p, input clk, output reg [7:0] mv);
    	integer state;
    	reg pe0_en,pe1_en,pe2_en,pe3_en,pe4_en,pe5_en,pe6_en,pe7_en,pe8_en,pe9_en,pe10_en,pe11_en,pe12_en,pe13_en,pe14_en,pe15_en;
    	reg [15:0] pe0_acc,pe1_acc,pe2_acc,pe3_acc,pe4_acc,pe5_acc,pe6_acc,pe7_acc,pe8_acc,pe9_acc,pe10_acc,pe11_acc,pe12_acc,pe13_acc,pe14_acc,pe15_acc;
	wire [7:0] pe0_out,pe1_out,pe2_out,pe3_out,pe4_out,pe5_out,pe6_out,pe7_out,pe8_out,pe9_out,pe10_out,pe11_out,pe12_out,pe13_out,pe14_out,pe15_out;

    	pe PE0(.a(c),.b(p),.en(pe0_en),.pe_out(pe0_out));
	pe PE1(.a(c),.b(p),.en(pe0_en),.pe_out(pe1_out));
	pe PE2(.a(c),.b(p),.en(pe0_en),.pe_out(pe2_out));
	pe PE3(.a(c),.b(p),.en(pe0_en),.pe_out(pe3_out));
	pe PE4(.a(c),.b(p),.en(pe0_en),.pe_out(pe4_out));
	pe PE5(.a(c),.b(p),.en(pe0_en),.pe_out(pe5_out));
	pe PE6(.a(c),.b(p),.en(pe0_en),.pe_out(pe6_out));
	pe PE7(.a(c),.b(p),.en(pe0_en),.pe_out(pe7_out));
	pe PE8(.a(c),.b(p),.en(pe0_en),.pe_out(pe8_out));
	pe PE9(.a(c),.b(p),.en(pe0_en),.pe_out(pe9_out));
	pe PE10(.a(c),.b(p),.en(pe0_en),.pe_out(pe10_out));
	pe PE11(.a(c),.b(p),.en(pe0_en),.pe_out(pe11_out));
	pe PE12(.a(c),.b(p),.en(pe0_en),.pe_out(pe12_out));
	pe PE13(.a(c),.b(p),.en(pe0_en),.pe_out(pe13_out));
	pe PE14(.a(c),.b(p),.en(pe0_en),.pe_out(pe14_out));
	pe PE15(.a(c),.b(p),.en(pe0_en),.pe_out(pe15_out));

	integer i;

    	initial begin
		pe0_acc = 16'd0;
		pe1_acc = 16'd0;
		pe2_acc = 16'd0;
		pe3_acc = 16'd0;
		pe4_acc = 16'd0;
		pe5_acc = 16'd0;
		pe6_acc = 16'd0;
		pe7_acc = 16'd0;
		pe8_acc = 16'd0;
		pe9_acc = 16'd0;
		pe10_acc = 16'd0;
		pe11_acc = 16'd0;
		pe12_acc = 16'd0;
		pe13_acc = 16'd0;
		pe14_acc = 16'd0;
		pe15_acc = 16'd0;
    	end
    	always @ (posedge clk) begin
        	for (i=0; i<272; i=i+1) begin
		state = i % 16;
		
		case (state)
            	0:  begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
                	state = 16;
			end
                	end
	    	1: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
			
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	2: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 1;
	       		state = 16;
			end
	       		end
	    	3: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end 
	    	4: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				state = 16;
			end
			else if (i >= 256) begin
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	5: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	6: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	7: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	8: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	9: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	10: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	11: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	12: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	13: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	14: begin
			if(i<16) begin
				pe0_en = 1;
				#50;
				pe0_acc = pe0_acc + pe0_out;
				pe1_en = 1;
				#50;
				pe1_acc = pe1_acc + pe1_out;
				pe2_en = 1;
				#50;
				pe2_acc = pe2_acc + pe2_out;
				pe3_en = 1;
				#50;
				pe3_acc = pe3_acc + pe3_out;
				pe4_en = 1;
				#50;
				pe4_acc = pe4_acc + pe4_out;
				$display("End of Sim: %d %d", i, pe4_out);
				pe5_en = 1;
				#50;
				pe5_acc = pe5_acc + pe5_out;
				pe6_en = 1;
				#50;
				pe6_acc = pe6_acc + pe6_out;
				pe7_en = 1;
				#50;
				pe7_acc = pe7_acc + pe7_out;
				pe8_en = 1;
				#50;
				pe8_acc = pe8_acc + pe8_out;
				pe9_en = 1;
				#50;
				pe9_acc = pe9_acc + pe9_out;
				pe10_en = 1;
				#50;
				pe10_acc = pe10_acc + pe10_out;
				pe11_en = 1;
				#50;
				pe11_acc = pe11_acc + pe11_out;
				pe12_en = 1;
				#50;
				pe12_acc = pe12_acc + pe12_out;
				pe13_en = 1;
				#50;
				pe13_acc = pe13_acc + pe13_out;
				pe14_en = 1;
				#50;
				pe14_acc = pe14_acc + pe14_out;
				state = 16;
			end
			else if (i >= 256) begin
				pe15_en = 1;
				#50;
				pe15_acc = pe15_acc + pe15_out;
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end
	    	15: begin
			if (i >= 256) begin
                		state = 16;
			end			
			else begin
			pe0_en = 1;
			#50;
			pe0_acc = pe0_acc + pe0_out;
			pe1_en = 1;
			#50;
			pe1_acc = pe1_acc + pe1_out;
			pe2_en = 1;
			#50;
			pe2_acc = pe2_acc + pe2_out;
			pe3_en = 1;
			#50;
			pe3_acc = pe3_acc + pe3_out;
			pe4_en = 1;
			#50;
			pe4_acc = pe4_acc + pe4_out;
			$display("End of Sim: %d %d", i, pe4_out);
			pe5_en = 1;
			#50;
			pe5_acc = pe5_acc + pe5_out;
			pe6_en = 1;
			#50;
			pe6_acc = pe6_acc + pe6_out;
			pe7_en = 1;
			#50;
			pe7_acc = pe7_acc + pe7_out;
			pe8_en = 1;
			#50;
			pe8_acc = pe8_acc + pe8_out;
			pe9_en = 1;
			#50;
			pe9_acc = pe9_acc + pe9_out;
			pe10_en = 1;
			#50;
			pe10_acc = pe10_acc + pe10_out;
			pe11_en = 1;
			#50;
			pe11_acc = pe11_acc + pe11_out;
			pe12_en = 1;
			#50;
			pe12_acc = pe12_acc + pe12_out;
			pe13_en = 1;
			#50;
			pe13_acc = pe13_acc + pe13_out;
			pe14_en = 1;
			#50;
			pe14_acc = pe14_acc + pe14_out;
			pe15_en = 1;
			#50;
			pe15_acc = pe15_acc + pe15_out;
	       		//pe0_en <= 0;
	       		state = 16;
			end
	       		end              
        	endcase
		end
    	end

	//assign mv = pe0_acc;

endmodule

module pe(input [7:0] a, input [7:0] b, input en, output reg [7:0] pe_out);
   	//reg [15:0] acc_temp = acc;
	always @* begin
	//$display("End of Sim: %d", en);
	if(en) begin
      		if (a<b) begin
        		assign pe_out = b - a;
      		end
      		else if (a==b) begin
        		assign pe_out = 8'd0;
      		end
      		else begin
        		assign pe_out = a - b;
      		end
		//acc_temp = acc_temp + pe_out;
		//acc = acc_temp;
		//$display("End of Sim: %d", acc);
	end
	else begin
		pe_out = 8'd0;	
	end
    	end
endmodule